// module mmio_dpi (
    
// );

// endmodule //mmio_dpi